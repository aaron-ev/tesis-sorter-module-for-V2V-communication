library verilog;
use verilog.vl_types.all;
entity smallSorter_vlg_vec_tst is
end smallSorter_vlg_vec_tst;
