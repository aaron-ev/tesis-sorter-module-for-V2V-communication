library verilog;
use verilog.vl_types.all;
entity trueDualPortRam_vlg_vec_tst is
end trueDualPortRam_vlg_vec_tst;
