library verilog;
use verilog.vl_types.all;
entity dist2Sorter_vlg_vec_tst is
end dist2Sorter_vlg_vec_tst;
