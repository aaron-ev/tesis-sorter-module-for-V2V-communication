library verilog;
use verilog.vl_types.all;
entity FSMDotProduct_vlg_vec_tst is
end FSMDotProduct_vlg_vec_tst;
