library verilog;
use verilog.vl_types.all;
entity dotProduct_vlg_vec_tst is
end dotProduct_vlg_vec_tst;
