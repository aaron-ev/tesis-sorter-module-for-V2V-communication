library verilog;
use verilog.vl_types.all;
entity merge8to16_vlg_vec_tst is
end merge8to16_vlg_vec_tst;
