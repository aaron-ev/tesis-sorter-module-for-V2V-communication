library verilog;
use verilog.vl_types.all;
entity dist2_vlg_vec_tst is
end dist2_vlg_vec_tst;
