

module complex2In4#(parameter WIDTH = 8)
(
	input clk, 
	input rst,
	input [WIDTH-1:0] inaReal,
	input [WIDTH-1:0] inaImag,
	input [WIDTH-1:0] inbReal,
	input [WIDTH-1:0] inbImag,
	input [WIDTH-1:0] incReal,
	input [WIDTH-1:0] incImag,	
	input [WIDTH-1:0] indReal,
	input [WIDTH-1:0] indImag,
	output [2*WIDTH-1:0] outaReal,
	output [2*WIDTH-1:0] outaImag,
	output [2*WIDTH-1:0] outbReal,
	output [2*WIDTH-1:0] outbImag,
	output [2*WIDTH-1:0] outcReal,
	output [2*WIDTH-1:0] outcImag,
	output [2*WIDTH-1:0] outdReal,
	output [2*WIDTH-1:0] outdImag	
);

complex2#(.WIDTH(8)) complex2a
(
	.clk(clk),
	.rst(rst),
	.aReal(inaReal),
	.aImag(inaImag),
	.outReal(outaReal),
	.outImag(outaImag)
);
complex2#(.WIDTH(8)) complex2b
(
	.clk(clk),
	.rst(rst),
	.aReal(inbReal),
	.aImag(inbImag),
	.outReal(outbReal),
	.outImag(outbImag)
);
complex2#(.WIDTH(8)) complex2c
(
	.clk(clk),
	.rst(rst),
	.aReal(incReal),
	.aImag(incImag),
	.outReal(outcReal),
	.outImag(outcImag)
);
complex2#(.WIDTH(8)) complex2d
(
	.clk(clk),
	.rst(rst),
	.aReal(indReal),
	.aImag(indImag),
	.outReal(outdReal),
	.outImag(outdImag)
);

endmodule