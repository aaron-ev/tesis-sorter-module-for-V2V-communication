library verilog;
use verilog.vl_types.all;
entity complexMul_vlg_vec_tst is
end complexMul_vlg_vec_tst;
