library verilog;
use verilog.vl_types.all;
entity merge4to8_vlg_vec_tst is
end merge4to8_vlg_vec_tst;
