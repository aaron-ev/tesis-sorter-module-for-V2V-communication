library verilog;
use verilog.vl_types.all;
entity regLoad_vlg_vec_tst is
end regLoad_vlg_vec_tst;
