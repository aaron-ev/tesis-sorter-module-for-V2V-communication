library verilog;
use verilog.vl_types.all;
entity complex2In4_vlg_vec_tst is
end complex2In4_vlg_vec_tst;
