library verilog;
use verilog.vl_types.all;
entity adderSub_vlg_vec_tst is
end adderSub_vlg_vec_tst;
