library verilog;
use verilog.vl_types.all;
entity m_2to4_vlg_vec_tst is
end m_2to4_vlg_vec_tst;
