library verilog;
use verilog.vl_types.all;
entity bufferTri_vlg_vec_tst is
end bufferTri_vlg_vec_tst;
