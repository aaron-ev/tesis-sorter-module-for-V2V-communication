library verilog;
use verilog.vl_types.all;
entity sortingNetwork4_vlg_vec_tst is
end sortingNetwork4_vlg_vec_tst;
