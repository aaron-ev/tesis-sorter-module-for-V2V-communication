library verilog;
use verilog.vl_types.all;
entity merge2to4_row_vlg_vec_tst is
end merge2to4_row_vlg_vec_tst;
