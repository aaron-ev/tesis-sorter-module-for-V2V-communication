library verilog;
use verilog.vl_types.all;
entity merge_vlg_vec_tst is
end merge_vlg_vec_tst;
