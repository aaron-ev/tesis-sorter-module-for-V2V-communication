library verilog;
use verilog.vl_types.all;
entity squareComplex_vlg_vec_tst is
end squareComplex_vlg_vec_tst;
