library verilog;
use verilog.vl_types.all;
entity ctrlUnitDotProduct_vlg_vec_tst is
end ctrlUnitDotProduct_vlg_vec_tst;
